../bexkat1/alu.sv