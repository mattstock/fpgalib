../bexkat1/intcalc.v