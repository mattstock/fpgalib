module registerfile
  #(WIDTH=32, COUNTP=4)
  (input              clk_i, 
   input 	      rst_i,
   input 	      supervisor, 
   input [COUNTP-1:0] read1,
   input [COUNTP-1:0] read2,
   input [COUNTP-1:0] write_addr,
   input [WIDTH-1:0]  write_data,
   input [1:0] 	      write_en,
   output [WIDTH-1:0] data1,
   output [WIDTH-1:0] data2);

  localparam COUNT=2**COUNTP;
  
  logic [WIDTH-1:0]   regfile [COUNT-1:0];
  logic [WIDTH-1:0]   regfile_next [COUNT-1:0];
  logic [WIDTH-1:0]   ssp, ssp_next;
  
  always_ff @(posedge clk_i or posedge rst_i)
    begin
      if (rst_i)
	begin
	  for (int i=0; i < COUNT; i = i + 1)
	    regfile[i] <= 'h00000000;
	  ssp <= 32'h0;
	end
      else
	begin
	  for (int i=0; i < COUNT; i = i + 1)
	    regfile[i] <= regfile_next[i];
	  ssp <= ssp_next;
	end // else: !if(rst_i)
    end // always_ff @

  always_comb
    begin
      for (int i=0; i < COUNT; i = i + 1)
	regfile_next[i] = regfile[i];
      ssp_next = ssp;
      data1 = (supervisor && read1 == 4'd15 ? ssp : regfile[read1]);
      data2 = (supervisor && read2 == 4'd15 ? ssp : regfile[read2]);
      case (write_en)
	2'b00: begin end
	2'b01:
	  begin
	    if (read1 == write_addr)
	      data1 = { 24'h0, write_data[7:0] };
	    if (read2 == write_addr)
	      data2 = { 24'h0, write_data[7:0] };
	    if (supervisor && write_addr == 4'd15)
	      ssp_next = { 24'h0, write_data[7:0] };
	    else
	      regfile_next[write_addr] = { 24'h000000, write_data[7:0] };
	  end
	2'b10:
	  begin
	    if (read1 == write_addr)
	      data1 = { 16'h0, write_data[15:0] };
	    if (read2 == write_addr)
	      data2 = { 16'h0, write_data[15:0] };
	    if (supervisor && write_addr == 4'd15)
	      ssp_next = { 16'h0, write_data[15:0] };
	    else
	      regfile_next[write_addr] = { 16'h0000, write_data[15:0] };
	  end
	2'b11:
	  begin
	    if (read1 == write_addr)
	      data1 = write_data;
	    if (read2 == write_addr)
	      data2 = write_data;
	    if (supervisor && write_addr == 4'd15)
	      ssp_next = write_data;
	    else
	      regfile_next[write_addr] = write_data;
	  end
      endcase // case (write_en)
    end // always_comb
endmodule // registerfile

