../bexkat1/alu.v