../../bexkat2/verilator/cache_top.sv